module hierarchy (input logic in1, in2, output logic out1, out2);
    comb c1(in1,in2,out1);
    comb c2(in1,in2,out2);
endmodule
